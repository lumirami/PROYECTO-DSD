// SISTEMA.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module SISTEMA (
		input  wire        clk_clk,                        
	   inout  				 scl,sda,
		input  wire        reset_reset_n,
		inout              HDMI_I2C_SCL,
      inout              HDMI_I2C_SDA,
      inout              HDMI_I2S,
      inout              HDMI_LRCLK,
      inout              HDMI_MCLK,
      inout              HDMI_SCLK,
      output             HDMI_TX_CLK,
      output      [23:0] HDMI_TX_D,
      output             HDMI_TX_DE,
      output             HDMI_TX_HS,
      input              HDMI_TX_INT,
      output             HDMI_TX_VS,
		input       [1:0]  KEY,
      output      [7:0]  LED 
	);

	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire  [19:0] cpu_data_master_address;                                   // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         cpu_data_master_read;                                      // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire         cpu_data_master_readdatavalid;                             // mm_interconnect_0:CPU_data_master_readdatavalid -> CPU:d_readdatavalid
	wire         cpu_data_master_write;                                     // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [31:0] cpu2_data_master_readdata;                                 // mm_interconnect_0:CPU2_data_master_readdata -> CPU2:d_readdata
	wire         cpu2_data_master_waitrequest;                              // mm_interconnect_0:CPU2_data_master_waitrequest -> CPU2:d_waitrequest
	wire         cpu2_data_master_debugaccess;                              // CPU2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU2_data_master_debugaccess
	wire  [19:0] cpu2_data_master_address;                                  // CPU2:d_address -> mm_interconnect_0:CPU2_data_master_address
	wire   [3:0] cpu2_data_master_byteenable;                               // CPU2:d_byteenable -> mm_interconnect_0:CPU2_data_master_byteenable
	wire         cpu2_data_master_read;                                     // CPU2:d_read -> mm_interconnect_0:CPU2_data_master_read
	wire         cpu2_data_master_write;                                    // CPU2:d_write -> mm_interconnect_0:CPU2_data_master_write
	wire  [31:0] cpu2_data_master_writedata;                                // CPU2:d_writedata -> mm_interconnect_0:CPU2_data_master_writedata
	wire  [31:0] cpu2_instruction_master_readdata;                          // mm_interconnect_0:CPU2_instruction_master_readdata -> CPU2:i_readdata
	wire         cpu2_instruction_master_waitrequest;                       // mm_interconnect_0:CPU2_instruction_master_waitrequest -> CPU2:i_waitrequest
	wire  [17:0] cpu2_instruction_master_address;                           // CPU2:i_address -> mm_interconnect_0:CPU2_instruction_master_address
	wire         cpu2_instruction_master_read;                              // CPU2:i_read -> mm_interconnect_0:CPU2_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [19:0] cpu_instruction_master_address;                            // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                               // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                      // mm_interconnect_0:CPU_instruction_master_readdatavalid -> CPU:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> JTAG_UART:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> JTAG_UART:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	wire  [31:0] mm_interconnect_0_sys_id_control_slave_readdata;           // SYS_ID:readdata -> mm_interconnect_0:SYS_ID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sys_id_control_slave_address;            // mm_interconnect_0:SYS_ID_control_slave_address -> SYS_ID:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                       // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                         // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [15:0] mm_interconnect_0_ram_s1_address;                          // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                       // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                            // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                        // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                            // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire  [31:0] mm_interconnect_0_data_counter_s1_readdata;                // data_counter:readdata -> mm_interconnect_0:data_counter_s1_readdata
	wire   [1:0] mm_interconnect_0_data_counter_s1_address;                 // mm_interconnect_0:data_counter_s1_address -> data_counter:address
	wire         mm_interconnect_0_share_m_s1_chipselect;                   // mm_interconnect_0:SHARE_M_s1_chipselect -> SHARE_M:chipselect
	wire  [31:0] mm_interconnect_0_share_m_s1_readdata;                     // SHARE_M:readdata -> mm_interconnect_0:SHARE_M_s1_readdata
	wire   [9:0] mm_interconnect_0_share_m_s1_address;                      // mm_interconnect_0:SHARE_M_s1_address -> SHARE_M:address
	wire   [3:0] mm_interconnect_0_share_m_s1_byteenable;                   // mm_interconnect_0:SHARE_M_s1_byteenable -> SHARE_M:byteenable
	wire         mm_interconnect_0_share_m_s1_write;                        // mm_interconnect_0:SHARE_M_s1_write -> SHARE_M:write
	wire  [31:0] mm_interconnect_0_share_m_s1_writedata;                    // mm_interconnect_0:SHARE_M_s1_writedata -> SHARE_M:writedata
	wire         mm_interconnect_0_share_m_s1_clken;                        // mm_interconnect_0:SHARE_M_s1_clken -> SHARE_M:clken
	wire         mm_interconnect_0_timer_0_s1_chipselect;                   // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                     // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                      // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                        // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                    // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire  [31:0] mm_interconnect_0_i2c_slave_s1_readdata;                   // i2c_slave:readdata -> mm_interconnect_0:i2c_slave_s1_readdata
	wire   [1:0] mm_interconnect_0_i2c_slave_s1_address;                    // mm_interconnect_0:i2c_slave_s1_address -> i2c_slave:address
	wire         mm_interconnect_0_hdmi_s1_chipselect;                      // mm_interconnect_0:HDMI_s1_chipselect -> HDMI:chipselect
	wire  [31:0] mm_interconnect_0_hdmi_s1_readdata;                        // HDMI:readdata -> mm_interconnect_0:HDMI_s1_readdata
	wire   [1:0] mm_interconnect_0_hdmi_s1_address;                         // mm_interconnect_0:HDMI_s1_address -> HDMI:address
	wire         mm_interconnect_0_hdmi_s1_write;                           // mm_interconnect_0:HDMI_s1_write -> HDMI:write_n
	wire  [31:0] mm_interconnect_0_hdmi_s1_writedata;                       // mm_interconnect_0:HDMI_s1_writedata -> HDMI:writedata
	wire  [31:0] mm_interconnect_0_cpu2_debug_mem_slave_readdata;           // CPU2:debug_mem_slave_readdata -> mm_interconnect_0:CPU2_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu2_debug_mem_slave_waitrequest;        // CPU2:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu2_debug_mem_slave_debugaccess;        // mm_interconnect_0:CPU2_debug_mem_slave_debugaccess -> CPU2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu2_debug_mem_slave_address;            // mm_interconnect_0:CPU2_debug_mem_slave_address -> CPU2:debug_mem_slave_address
	wire         mm_interconnect_0_cpu2_debug_mem_slave_read;               // mm_interconnect_0:CPU2_debug_mem_slave_read -> CPU2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu2_debug_mem_slave_byteenable;         // mm_interconnect_0:CPU2_debug_mem_slave_byteenable -> CPU2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu2_debug_mem_slave_write;              // mm_interconnect_0:CPU2_debug_mem_slave_write -> CPU2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu2_debug_mem_slave_writedata;          // mm_interconnect_0:CPU2_debug_mem_slave_writedata -> CPU2:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram2_s1_chipselect;                      // mm_interconnect_0:RAM2_s1_chipselect -> RAM2:chipselect
	wire  [31:0] mm_interconnect_0_ram2_s1_readdata;                        // RAM2:readdata -> mm_interconnect_0:RAM2_s1_readdata
	wire  [13:0] mm_interconnect_0_ram2_s1_address;                         // mm_interconnect_0:RAM2_s1_address -> RAM2:address
	wire   [3:0] mm_interconnect_0_ram2_s1_byteenable;                      // mm_interconnect_0:RAM2_s1_byteenable -> RAM2:byteenable
	wire         mm_interconnect_0_ram2_s1_write;                           // mm_interconnect_0:RAM2_s1_write -> RAM2:write
	wire  [31:0] mm_interconnect_0_ram2_s1_writedata;                       // mm_interconnect_0:RAM2_s1_writedata -> RAM2:writedata
	wire         mm_interconnect_0_ram2_s1_clken;                           // mm_interconnect_0:RAM2_s1_clken -> RAM2:clken
	wire         mm_interconnect_0_share_m_s2_chipselect;                   // mm_interconnect_0:SHARE_M_s2_chipselect -> SHARE_M:chipselect2
	wire  [31:0] mm_interconnect_0_share_m_s2_readdata;                     // SHARE_M:readdata2 -> mm_interconnect_0:SHARE_M_s2_readdata
	wire   [9:0] mm_interconnect_0_share_m_s2_address;                      // mm_interconnect_0:SHARE_M_s2_address -> SHARE_M:address2
	wire   [3:0] mm_interconnect_0_share_m_s2_byteenable;                   // mm_interconnect_0:SHARE_M_s2_byteenable -> SHARE_M:byteenable2
	wire         mm_interconnect_0_share_m_s2_write;                        // mm_interconnect_0:SHARE_M_s2_write -> SHARE_M:write2
	wire  [31:0] mm_interconnect_0_share_m_s2_writedata;                    // mm_interconnect_0:SHARE_M_s2_writedata -> SHARE_M:writedata2
	wire         mm_interconnect_0_share_m_s2_clken;                        // mm_interconnect_0:SHARE_M_s2_clken -> SHARE_M:clken2
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> CPU:irq
	wire  [31:0] cpu2_irq_irq;                                              // irq_mapper_001:sender_irq -> CPU2:irq
	wire         irq_mapper_receiver0_irq;                                  // JTAG_UART:av_irq -> [irq_mapper:receiver0_irq, irq_mapper_001:receiver0_irq]
	wire         irq_mapper_receiver1_irq;                                  // timer_0:irq -> [irq_mapper:receiver1_irq, irq_mapper_001:receiver1_irq]
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [CPU:reset_n, irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [CPU:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                             // CPU:debug_reset_request -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [CPU2:reset_n, irq_mapper_001:reset, mm_interconnect_0:CPU2_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset_req;                    // rst_controller_001:reset_req -> [CPU2:reset_req, rst_translator_001:reset_req_in]
	wire         cpu2_debug_reset_request_reset;                            // CPU2:debug_reset_request -> rst_controller_001:reset_in1
	wire         rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [HDMI:reset_n, JTAG_UART:rst_n, RAM2:reset, RAM:reset, SHARE_M:reset, SYS_ID:reset_n, data_counter:reset_n, i2c_slave:reset_n, mm_interconnect_0:JTAG_UART_reset_reset_bridge_in_reset_reset, rst_translator_002:in_reset, timer_0:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                    // rst_controller_002:reset_req -> [RAM2:reset_req, RAM:reset_req, SHARE_M:reset_req, rst_translator_002:reset_req_in]
	wire			 c_up;
	wire [12:0]  data_counter_external_connection_export;
	wire [7:0]   i2c_slave_export;
	wire [2:0]   selector_export;
	SISTEMA_CPU cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	SISTEMA_CPU2 cpu2 (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),             //                          .reset_req
		.d_address                           (cpu2_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu2_data_master_read),                              //                          .read
		.d_readdata                          (cpu2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu2_data_master_write),                             //                          .write
		.d_writedata                         (cpu2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu2_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	SISTEMA_HDMI hdmi (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_hdmi_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hdmi_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hdmi_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hdmi_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hdmi_s1_readdata),   //                    .readdata
		.out_port   (selector_export)                       // external_connection.export
	);

	SISTEMA_JTAG_UART jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	SISTEMA_RAM ram (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),       //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),         //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect),    //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),         //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),      //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),     //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable),    //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req), //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	SISTEMA_RAM2 ram2 (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_ram2_s1_address),      //     s1.address
		.clken      (mm_interconnect_0_ram2_s1_clken),        //       .clken
		.chipselect (mm_interconnect_0_ram2_s1_chipselect),   //       .chipselect
		.write      (mm_interconnect_0_ram2_s1_write),        //       .write
		.readdata   (mm_interconnect_0_ram2_s1_readdata),     //       .readdata
		.writedata  (mm_interconnect_0_ram2_s1_writedata),    //       .writedata
		.byteenable (mm_interconnect_0_ram2_s1_byteenable),   //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req), //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	SISTEMA_SHARE_M share_m (
		.address     (mm_interconnect_0_share_m_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_share_m_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_share_m_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_share_m_s1_write),      //       .write
		.readdata    (mm_interconnect_0_share_m_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_share_m_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_share_m_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_0_share_m_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_share_m_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_share_m_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_share_m_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_share_m_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_share_m_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_share_m_s2_byteenable), //       .byteenable
		.clk         (clk_clk),                                 //   clk1.clk
		.reset       (rst_controller_002_reset_out_reset),      // reset1.reset
		.reset_req   (rst_controller_002_reset_out_reset_req),  //       .reset_req
		.freeze      (1'b0)                                     // (terminated)
	);

	SISTEMA_SYS_ID sys_id (
		.clock    (clk_clk),                                         //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),             //         reset.reset_n
		.readdata (mm_interconnect_0_sys_id_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sys_id_control_slave_address)   //              .address
	);
counter				 u_counter		 (
		.up(c_up),
		.nrst(reset_reset_n),
		.q(data_counter_external_connection_export)
	);
I2C_slave				u_I2C_slave(
		.scl(scl),
		.sda(sda),
		.clk(clk_clk),
		.rst(reset_reset_n),
		.data_valid(c_up),
		.data_from_master(i2c_slave_export)
	);
DE10_Nano_HDMI_TX		u_HDMI		(
	   .FPGA_CLK1_50(clk_clk),
      .HDMI_I2C_SCL(HDMI_I2C_SCL),
      .HDMI_I2C_SDA(HDMI_I2C_SDA),
      .HDMI_I2S(HDMI_I2S),
      .HDMI_LRCLK(HDMI_LRCLK),
      .HDMI_MCLK(HDMI_MCLK),
      .HDMI_SCLK(HDMI_SCLK),
      .HDMI_TX_CLK(HDMI_TX_CLK),
      .HDMI_TX_D(HDMI_TX_D),
      .HDMI_TX_DE(HDMI_TX_DE),
      .HDMI_TX_HS(HDMI_TX_HS),
      .HDMI_TX_INT(HDMI_TX_INT),
      .HDMI_TX_VS(HDMI_TX_VS),
      .KEY(KEY),
      .LED(LED),
      .SW(selector_export)
	);
	SISTEMA_data_counter data_counter (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_data_counter_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_data_counter_s1_readdata), //                    .readdata
		.in_port  (data_counter_external_connection_export)     // external_connection.export
	);

	SISTEMA_i2c_slave i2c_slave (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_i2c_slave_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_i2c_slave_s1_readdata), //                    .readdata
		.in_port  (i2c_slave_export)                         // external_connection.export
	);

	SISTEMA_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	SISTEMA_mm_interconnect_0 mm_interconnect_0 (
		.CLK_50_clk_clk                              (clk_clk),                                                   //                            CLK_50_clk.clk
		.CPU2_reset_reset_bridge_in_reset_reset      (rst_controller_001_reset_out_reset),                        //      CPU2_reset_reset_bridge_in_reset.reset
		.CPU_reset_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                            //       CPU_reset_reset_bridge_in_reset.reset
		.JTAG_UART_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                        // JTAG_UART_reset_reset_bridge_in_reset.reset
		.CPU_data_master_address                     (cpu_data_master_address),                                   //                       CPU_data_master.address
		.CPU_data_master_waitrequest                 (cpu_data_master_waitrequest),                               //                                      .waitrequest
		.CPU_data_master_byteenable                  (cpu_data_master_byteenable),                                //                                      .byteenable
		.CPU_data_master_read                        (cpu_data_master_read),                                      //                                      .read
		.CPU_data_master_readdata                    (cpu_data_master_readdata),                                  //                                      .readdata
		.CPU_data_master_readdatavalid               (cpu_data_master_readdatavalid),                             //                                      .readdatavalid
		.CPU_data_master_write                       (cpu_data_master_write),                                     //                                      .write
		.CPU_data_master_writedata                   (cpu_data_master_writedata),                                 //                                      .writedata
		.CPU_data_master_debugaccess                 (cpu_data_master_debugaccess),                               //                                      .debugaccess
		.CPU_instruction_master_address              (cpu_instruction_master_address),                            //                CPU_instruction_master.address
		.CPU_instruction_master_waitrequest          (cpu_instruction_master_waitrequest),                        //                                      .waitrequest
		.CPU_instruction_master_read                 (cpu_instruction_master_read),                               //                                      .read
		.CPU_instruction_master_readdata             (cpu_instruction_master_readdata),                           //                                      .readdata
		.CPU_instruction_master_readdatavalid        (cpu_instruction_master_readdatavalid),                      //                                      .readdatavalid
		.CPU2_data_master_address                    (cpu2_data_master_address),                                  //                      CPU2_data_master.address
		.CPU2_data_master_waitrequest                (cpu2_data_master_waitrequest),                              //                                      .waitrequest
		.CPU2_data_master_byteenable                 (cpu2_data_master_byteenable),                               //                                      .byteenable
		.CPU2_data_master_read                       (cpu2_data_master_read),                                     //                                      .read
		.CPU2_data_master_readdata                   (cpu2_data_master_readdata),                                 //                                      .readdata
		.CPU2_data_master_write                      (cpu2_data_master_write),                                    //                                      .write
		.CPU2_data_master_writedata                  (cpu2_data_master_writedata),                                //                                      .writedata
		.CPU2_data_master_debugaccess                (cpu2_data_master_debugaccess),                              //                                      .debugaccess
		.CPU2_instruction_master_address             (cpu2_instruction_master_address),                           //               CPU2_instruction_master.address
		.CPU2_instruction_master_waitrequest         (cpu2_instruction_master_waitrequest),                       //                                      .waitrequest
		.CPU2_instruction_master_read                (cpu2_instruction_master_read),                              //                                      .read
		.CPU2_instruction_master_readdata            (cpu2_instruction_master_readdata),                          //                                      .readdata
		.CPU_debug_mem_slave_address                 (mm_interconnect_0_cpu_debug_mem_slave_address),             //                   CPU_debug_mem_slave.address
		.CPU_debug_mem_slave_write                   (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                      .write
		.CPU_debug_mem_slave_read                    (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                      .read
		.CPU_debug_mem_slave_readdata                (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                      .readdata
		.CPU_debug_mem_slave_writedata               (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                      .writedata
		.CPU_debug_mem_slave_byteenable              (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                      .byteenable
		.CPU_debug_mem_slave_waitrequest             (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                      .waitrequest
		.CPU_debug_mem_slave_debugaccess             (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                      .debugaccess
		.CPU2_debug_mem_slave_address                (mm_interconnect_0_cpu2_debug_mem_slave_address),            //                  CPU2_debug_mem_slave.address
		.CPU2_debug_mem_slave_write                  (mm_interconnect_0_cpu2_debug_mem_slave_write),              //                                      .write
		.CPU2_debug_mem_slave_read                   (mm_interconnect_0_cpu2_debug_mem_slave_read),               //                                      .read
		.CPU2_debug_mem_slave_readdata               (mm_interconnect_0_cpu2_debug_mem_slave_readdata),           //                                      .readdata
		.CPU2_debug_mem_slave_writedata              (mm_interconnect_0_cpu2_debug_mem_slave_writedata),          //                                      .writedata
		.CPU2_debug_mem_slave_byteenable             (mm_interconnect_0_cpu2_debug_mem_slave_byteenable),         //                                      .byteenable
		.CPU2_debug_mem_slave_waitrequest            (mm_interconnect_0_cpu2_debug_mem_slave_waitrequest),        //                                      .waitrequest
		.CPU2_debug_mem_slave_debugaccess            (mm_interconnect_0_cpu2_debug_mem_slave_debugaccess),        //                                      .debugaccess
		.data_counter_s1_address                     (mm_interconnect_0_data_counter_s1_address),                 //                       data_counter_s1.address
		.data_counter_s1_readdata                    (mm_interconnect_0_data_counter_s1_readdata),                //                                      .readdata
		.HDMI_s1_address                             (mm_interconnect_0_hdmi_s1_address),                         //                               HDMI_s1.address
		.HDMI_s1_write                               (mm_interconnect_0_hdmi_s1_write),                           //                                      .write
		.HDMI_s1_readdata                            (mm_interconnect_0_hdmi_s1_readdata),                        //                                      .readdata
		.HDMI_s1_writedata                           (mm_interconnect_0_hdmi_s1_writedata),                       //                                      .writedata
		.HDMI_s1_chipselect                          (mm_interconnect_0_hdmi_s1_chipselect),                      //                                      .chipselect
		.i2c_slave_s1_address                        (mm_interconnect_0_i2c_slave_s1_address),                    //                          i2c_slave_s1.address
		.i2c_slave_s1_readdata                       (mm_interconnect_0_i2c_slave_s1_readdata),                   //                                      .readdata
		.JTAG_UART_avalon_jtag_slave_address         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //           JTAG_UART_avalon_jtag_slave.address
		.JTAG_UART_avalon_jtag_slave_write           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                      .write
		.JTAG_UART_avalon_jtag_slave_read            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                      .read
		.JTAG_UART_avalon_jtag_slave_readdata        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                      .readdata
		.JTAG_UART_avalon_jtag_slave_writedata       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                      .writedata
		.JTAG_UART_avalon_jtag_slave_waitrequest     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                      .waitrequest
		.JTAG_UART_avalon_jtag_slave_chipselect      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                      .chipselect
		.RAM_s1_address                              (mm_interconnect_0_ram_s1_address),                          //                                RAM_s1.address
		.RAM_s1_write                                (mm_interconnect_0_ram_s1_write),                            //                                      .write
		.RAM_s1_readdata                             (mm_interconnect_0_ram_s1_readdata),                         //                                      .readdata
		.RAM_s1_writedata                            (mm_interconnect_0_ram_s1_writedata),                        //                                      .writedata
		.RAM_s1_byteenable                           (mm_interconnect_0_ram_s1_byteenable),                       //                                      .byteenable
		.RAM_s1_chipselect                           (mm_interconnect_0_ram_s1_chipselect),                       //                                      .chipselect
		.RAM_s1_clken                                (mm_interconnect_0_ram_s1_clken),                            //                                      .clken
		.RAM2_s1_address                             (mm_interconnect_0_ram2_s1_address),                         //                               RAM2_s1.address
		.RAM2_s1_write                               (mm_interconnect_0_ram2_s1_write),                           //                                      .write
		.RAM2_s1_readdata                            (mm_interconnect_0_ram2_s1_readdata),                        //                                      .readdata
		.RAM2_s1_writedata                           (mm_interconnect_0_ram2_s1_writedata),                       //                                      .writedata
		.RAM2_s1_byteenable                          (mm_interconnect_0_ram2_s1_byteenable),                      //                                      .byteenable
		.RAM2_s1_chipselect                          (mm_interconnect_0_ram2_s1_chipselect),                      //                                      .chipselect
		.RAM2_s1_clken                               (mm_interconnect_0_ram2_s1_clken),                           //                                      .clken
		.SHARE_M_s1_address                          (mm_interconnect_0_share_m_s1_address),                      //                            SHARE_M_s1.address
		.SHARE_M_s1_write                            (mm_interconnect_0_share_m_s1_write),                        //                                      .write
		.SHARE_M_s1_readdata                         (mm_interconnect_0_share_m_s1_readdata),                     //                                      .readdata
		.SHARE_M_s1_writedata                        (mm_interconnect_0_share_m_s1_writedata),                    //                                      .writedata
		.SHARE_M_s1_byteenable                       (mm_interconnect_0_share_m_s1_byteenable),                   //                                      .byteenable
		.SHARE_M_s1_chipselect                       (mm_interconnect_0_share_m_s1_chipselect),                   //                                      .chipselect
		.SHARE_M_s1_clken                            (mm_interconnect_0_share_m_s1_clken),                        //                                      .clken
		.SHARE_M_s2_address                          (mm_interconnect_0_share_m_s2_address),                      //                            SHARE_M_s2.address
		.SHARE_M_s2_write                            (mm_interconnect_0_share_m_s2_write),                        //                                      .write
		.SHARE_M_s2_readdata                         (mm_interconnect_0_share_m_s2_readdata),                     //                                      .readdata
		.SHARE_M_s2_writedata                        (mm_interconnect_0_share_m_s2_writedata),                    //                                      .writedata
		.SHARE_M_s2_byteenable                       (mm_interconnect_0_share_m_s2_byteenable),                   //                                      .byteenable
		.SHARE_M_s2_chipselect                       (mm_interconnect_0_share_m_s2_chipselect),                   //                                      .chipselect
		.SHARE_M_s2_clken                            (mm_interconnect_0_share_m_s2_clken),                        //                                      .clken
		.SYS_ID_control_slave_address                (mm_interconnect_0_sys_id_control_slave_address),            //                  SYS_ID_control_slave.address
		.SYS_ID_control_slave_readdata               (mm_interconnect_0_sys_id_control_slave_readdata),           //                                      .readdata
		.timer_0_s1_address                          (mm_interconnect_0_timer_0_s1_address),                      //                            timer_0_s1.address
		.timer_0_s1_write                            (mm_interconnect_0_timer_0_s1_write),                        //                                      .write
		.timer_0_s1_readdata                         (mm_interconnect_0_timer_0_s1_readdata),                     //                                      .readdata
		.timer_0_s1_writedata                        (mm_interconnect_0_timer_0_s1_writedata),                    //                                      .writedata
		.timer_0_s1_chipselect                       (mm_interconnect_0_timer_0_s1_chipselect)                    //                                      .chipselect
	);

	SISTEMA_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	SISTEMA_irq_mapper irq_mapper_001 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (cpu2_irq_irq)                        //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu2_debug_reset_request_reset),         // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
